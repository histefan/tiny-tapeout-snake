module draw_snake #(
    parameter SIZE = 5,
    parameter BIT = 10,
    parameter X_START = 320, // start position of snake
    parameter Y_START = 240
) (
    input wire clk,
    input wire reset,
    input wire update,
    input wire[BIT-1:0] x_pos,
    input wire[BIT-1:0] y_pos, 
    input wire [2:0] direction,
    input wire [1:0] game_state,  
    output wire snake_head_active,
    output wire snake_body_active,
    output wire [2:0] rgb
);

parameter snake_rgb = 3'b010; // green


// states control
localparam IDLE = 3'b000;
localparam UP = 3'b001;
localparam DOWN = 3'b010;
localparam LEFT = 3'b011;
localparam RIGHT = 3'b100;

//states game
localparam PLAY = 2'b01;
localparam GAME_OVER = 2'b11;

integer i,j;
reg [BIT-1:0] snakeX, next_snakeX, snakeY, next_snakeY; 
reg [BIT-1:0] bodyX [0:31];
reg [BIT-1:0] bodyY [0:31];
reg [BIT-1:0] next_bodyX [0:31];
reg [BIT-1:0] next_bodyY [0:31];  //, next_bodyX1, next_bodyX2;

always @(posedge clk) begin
    if (reset) begin
        //size <= 5'b00001;
        snakeX <= X_START;
        snakeY <= Y_START;
         for (i = 0; i < 32; i = i+1) begin
            bodyX[i] <= 10'd700;
            bodyY[i] <= 10'd500;   
        end        
    end else begin
        snakeX <= next_snakeX;
        snakeY <= next_snakeY;
        for (i = 0; i < 32; i = i+1) begin
            bodyX[i] <= next_bodyX[i];
            bodyY[i] <= next_bodyY[i];   
        end
        //size <= next_size;
    end
end

always @(snakeX, snakeY, game_state, direction, update, bodyX[0], bodyY[0]) begin
    next_snakeX = snakeX;
    next_snakeY = snakeY;
    for (i = 0; i < 32; i = i+1) begin
            next_bodyX[i] = bodyX[i];
            next_bodyY[i] = bodyY[i];   
    end
    
    //next_size = size;
    if (game_state == PLAY && update) begin
            // shift values in register
            case (direction) // direction of head
            UP: next_snakeY = (snakeY - SIZE);
            DOWN: next_snakeY = (snakeY + SIZE);
            LEFT : next_snakeX = (snakeX - SIZE);
            RIGHT: next_snakeX = (snakeX + SIZE);
            IDLE: begin 
                    next_snakeY = snakeY;
                    next_snakeX = snakeX;
                  end
            default:begin 
                    next_snakeY = snakeY;
                    next_snakeX = snakeX;
                  end
        endcase 
        for (j = 1; j < 32; j = j+1) begin
            next_bodyX[j] = bodyX[j-1];
            next_bodyY[j] = bodyY[j-1];   
        end
        next_bodyX[0] = snakeX;
        next_bodyY[0] = snakeY;
        
    end     
    if (game_state == GAME_OVER)  begin  
        //initialise snake head
        //next_size = 5'b00010;
        next_snakeX = X_START;
        next_snakeY = Y_START;    
    end    
end

assign snake_head_active = (x_pos >= snakeX) && (x_pos < snakeX + SIZE) && (y_pos >= snakeY) && (y_pos < snakeY + SIZE);
//assign snake_head_active = (x_pos >= snakeX) && (x_pos < snakeX + SIZE) && (y_pos >= snakeY) && (y_pos < snakeY + SIZE);


//temporary
assign snake_body_active = (x_pos >= bodyX[0]) && (x_pos < bodyX[0] + SIZE) && (y_pos >= bodyY[0]) && (y_pos < bodyY[0] + SIZE) ||
(x_pos >= bodyX[1]) && (x_pos < bodyX[1] + SIZE) && (y_pos >= bodyY[1]) && (y_pos < bodyY[1] + SIZE) ||
(x_pos >= bodyX[2]) && (x_pos < bodyX[2] + SIZE) && (y_pos >= bodyY[2]) && (y_pos < bodyY[2] + SIZE) ||
(x_pos >= bodyX[3]) && (x_pos < bodyX[3] + SIZE) && (y_pos >= bodyY[3]) && (y_pos < bodyY[3] + SIZE) ||
(x_pos >= bodyX[4]) && (x_pos < bodyX[4] + SIZE) && (y_pos >= bodyY[4]) && (y_pos < bodyY[4] + SIZE);


assign rgb = snake_rgb;




 
endmodule
